class eth_packet_sw extends uvm_sequence_item;

endclass : eth_packet_sw