class configuration extends uvm_object;
    virtual eth_if_in.inp vif_in;
    `uvm_object_utils(configuration)
    
endclass : configuration